module color(clk, rst, q);
   input clk;
   input rst;
   output [7:0] q;
   reg [7:0]    q;
   reg [5:0]    s;
   
   always @(posedge clk or negedge rst)
      if (!rst)
         s <= 6'b000000;
      else if(clk==1)
      begin
         if (s == 6'b101101)
            s <= 6'b000000;
         else
			begin
            s <= s + 6'b000001;
         case (s)
      ///////////第一种花形
				6'b000000 :
               q <= 8'b00000000;
					
            6'b000001 :
               q <= 8'b10000001;
            6'b000010 :
               q <= 8'b01000010;
            6'b000011 :
               q <= 8'b00100100;
            6'b000100 :
               q <= 8'b00011000;
            6'b000101 :
               q <= 8'b00000000;
		///////////第二种花形
            6'b000110 :
               q <= 8'b00011000;
            6'b000111 :
               q <= 8'b00111100;
            6'b001000 :
               q <= 8'b01111110;
            6'b001001 :
               q <= 8'b11111111;
            6'b001010 :
               q <= 8'b11100111;
            6'b001011 :
               q <= 8'b11000011;
            6'b001100 :
               q <= 8'b10000001;
            6'b001101 :
               q <= 8'b00000000;
		///////////第三种花型
            6'b001110 :
               q <= 8'b10000000;
            6'b001111 :
               q <= 8'b11000000;
            6'b010000 :
               q <= 8'b11100000;
            6'b010001 :
               q <= 8'b11110000;
            6'b010010 :
               q <= 8'b11111000;
            6'b010011 :
               q <= 8'b11111100;
            6'b010100 :
               q <= 8'b11111110;
            6'b010101 :
               q <= 8'b11111111;
            6'b010110 :
               q <= 8'b11111110;
            6'b010111 :
               q <= 8'b11111100;
            6'b011000 :
               q <= 8'b11111000;
            6'b011001 :
               q <= 8'b11110000;
            6'b011010 :
               q <= 8'b11100000;
            6'b011011 :
               q <= 8'b11000000;
            6'b011100 :
               q <= 8'b10000000;
            6'b011101 :
               q <= 8'b00000000;
		///////////第四种花型
				6'b011110 :
               q <= 8'b00000001;
            6'b011111 :
               q <= 8'b00000011;
            6'b100000 :
               q <= 8'b00000111;
            6'b100001 :
               q <= 8'b00001111;
            6'b100010 :
               q <= 8'b00011111;
            6'b100011 :
               q <= 8'b00111111;
            6'b100100 :
               q <= 8'b01111111;
            6'b100101 :
               q <= 8'b11111111;
            6'b100110 :
               q <= 8'b01111111;
            6'b100111 :
               q <= 8'b00111111;
            6'b101000 :
               q <= 8'b00011111;
            6'b101001 :
               q <= 8'b00001111;
            6'b101010 :
               q <= 8'b00000111;
            6'b101011 :
               q <= 8'b00000011;
            6'b101100 :
               q <= 8'b00000001;
            6'b101101 :
               q <= 8'b00000000;
            default :
               ;
         endcase
			end
      end
   
endmodule
